module Player (
input nrst,
input clk,
output reg	map_counter,
output reg	time_counter,
output reg	eight_note
);


always @( posedge clk or negedge nrst) begin
	
end

endmodule